module tamrin_1(input a,b,c,d,e,output y,z);
    assign y= ~c;
    assign z=(a&b);
endmodule
