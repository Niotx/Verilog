`timescale 1ns/100ps
module Q4_TB();
    reg X1,X2,X3,X4,X5;
    wire FFINAL , GFINAL;
    Q4_1 testf(.x1(X1),.x2(X2),.x3(X3),.x4(X4),.x5(X5),.ffinal(FFINAL));
    Q4_2 testg(.x1(X1),.x2(X2),.x3(X3),.x4(X4),.x5(X5),.gfinal(GFINAL));
    initial begin 
        X1 <= 0 ; X2 <= 0 ;
        X3 <= 0 ; X4 <= 0 ;
        X5 <= 0 ;

        #100

        X1 <= 0 ; X2 <= 0 ;
        X3 <= 0 ; X4 <= 0 ;
        X5 <= 1 ;

        #100

        X1 <= 0 ; X2 <= 0 ;
        X3 <= 0 ; X4 <= 1 ;
        X5 <= 0 ;

        #100

        X1 <= 0 ; X2 <= 0 ;
        X3 <= 0 ; X4 <= 1 ;
        X5 <= 1 ;

        #100

        X1 <= 0 ; X2 <= 0 ;
        X3 <= 1 ; X4 <= 0 ;
        X5 <= 0 ;

        #100

        X1 <= 0 ; X2 <= 0 ;
        X3 <= 1 ; X4 <= 0 ;
        X5 <= 1 ;

        #100

        X1 <= 0 ; X2 <= 0 ;
        X3 <= 1 ; X4 <= 1 ;
        X5 <= 0 ;

        #100

        X1 <= 0 ; X2 <= 0 ;
        X3 <= 1 ; X4 <= 1 ;
        X5 <= 1 ;

        #100

        X1 <= 0 ; X2 <= 1 ;
        X3 <= 0 ; X4 <= 0 ;
        X5 <= 0 ;

        #100

        X1 <= 0 ; X2 <= 1 ;
        X3 <= 0 ; X4 <= 0 ;
        X5 <= 1 ;

        #100

        X1 <= 0 ; X2 <= 1 ;
        X3 <= 0 ; X4 <= 1 ;
        X5 <= 0 ;

        #100

        X1 <= 0 ; X2 <= 1 ;
        X3 <= 0 ; X4 <= 1 ;
        X5 <= 1 ;

        #100

        X1 <= 0 ; X2 <= 1 ;
        X3 <= 1 ; X4 <= 0 ;
        X5 <= 0 ;

        #100

        X1 <= 0 ; X2 <= 1 ;
        X3 <= 1 ; X4 <= 0 ;
        X5 <= 1 ;

        #100

        X1 <= 0 ; X2 <= 1 ;
        X3 <= 1 ; X4 <= 1 ;
        X5 <= 0 ;

        #100

        X1 <= 0 ; X2 <= 1 ;
        X3 <= 1 ; X4 <= 1 ;
        X5 <= 1 ;

        #100

        X1 <= 1 ; X2 <= 0 ;
        X3 <= 0 ; X4 <= 0 ;
        X5 <= 0 ;

        #100

        X1 <= 1 ; X2 <= 0 ;
        X3 <= 0 ; X4 <= 0 ;
        X5 <= 1 ;

        #100

        X1 <= 1 ; X2 <= 0 ;
        X3 <= 0 ; X4 <= 1 ;
        X5 <= 0 ;

        #100

        X1 <= 1 ; X2 <= 0 ;
        X3 <= 0 ; X4 <= 1 ;
        X5 <= 1 ;

        #100

        X1 <= 1 ; X2 <= 0 ;
        X3 <= 1 ; X4 <= 0 ;
        X5 <= 0 ;

        #100

        X1 <= 1 ; X2 <= 0 ;
        X3 <= 1 ; X4 <= 0 ;
        X5 <= 1 ;

        #100

        X1 <= 1 ; X2 <= 0 ;
        X3 <= 1 ; X4 <= 1 ;
        X5 <= 0 ;

        #100

        X1 <= 1 ; X2 <= 0 ;
        X3 <= 1 ; X4 <= 1 ;
        X5 <= 1 ;

        #100

        X1 <= 1 ; X2 <= 1 ;
        X3 <= 0 ; X4 <= 0 ;
        X5 <= 0 ;

        #100

        X1 <= 1 ; X2 <= 1 ;
        X3 <= 0 ; X4 <= 0 ;
        X5 <= 1 ;

        #100

        X1 <= 1 ; X2 <= 1 ;
        X3 <= 0 ; X4 <= 1 ;
        X5 <= 0 ;

        #100

        X1 <= 1 ; X2 <= 1 ;
        X3 <= 0 ; X4 <= 1 ;
        X5 <= 1 ;

        #100

        X1 <= 1 ; X2 <= 1 ;
        X3 <= 1 ; X4 <= 0 ;
        X5 <= 0 ;

        #100

        X1 <= 1 ; X2 <= 1 ;
        X3 <= 1 ; X4 <= 0 ;
        X5 <= 1 ;

        #100

        X1 <= 1 ; X2 <= 1 ;
        X3 <= 1 ; X4 <= 1 ;
        X5 <= 0 ;

        #100

        X1 <= 1 ; X2 <= 1 ;
        X3 <= 1 ; X4 <= 1 ;
        X5 <= 1 ;

        #100;
    end
endmodule